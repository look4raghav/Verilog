module test (input [7:0] a,
						 b,
			 output [7:0] c);
endmodule

module test ( input wire [7:0] a,
			  input wire [7:0] b,
			  output reg [7:0] c);
endmodule