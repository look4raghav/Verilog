module <name> ([port_list]);
  
endmodule

module name;
  
endmodule