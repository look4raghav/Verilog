module (input a,
				b,
		output c);

endmodule


module ( input signed a, b,
         output c);
    wire a, b;
    reg signed c;
endmodule;