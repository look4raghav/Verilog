module my_design (input wire clk,
				  input en,
				  input rw,
				  input [15:0] data,
				  output int);

endmodule