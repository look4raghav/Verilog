module tb;
  initial
    $display("Hello World !");
  endmodule