module testbench;
  design d0 ( [port_list_connections] );
endmodule